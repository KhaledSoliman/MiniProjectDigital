module timer (S_ADR_I, S_DAT_I, S_WE_I, S_STB_I, S_CYC_I, S_CTI_I, S_BTE_I, S_LOCK_I, S_SEL_I, CLK_I, RST_I, S_DAT_O, S_ACK_O, S_RTY_O, S_ERR_O, S_INT_O, RSTREQ_O, TOPULSE_O);

input S_WE_I;
input S_STB_I;
input S_CYC_I;
input S_LOCK_I;
input CLK_I;
input RST_I;
output S_ACK_O;
output S_RTY_O;
output S_ERR_O;
output S_INT_O;
output RSTREQ_O;
output TOPULSE_O;
input [31:0] S_ADR_I;
input [31:0] S_DAT_I;
input [2:0] S_CTI_I;
input [1:0] S_BTE_I;
input [3:0] S_SEL_I;
output [31:0] S_DAT_O;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX4 BUFX4_1 ( .A(_13_), .Y(_13__bF_buf4) );
BUFX4 BUFX4_2 ( .A(_13_), .Y(_13__bF_buf3) );
BUFX4 BUFX4_3 ( .A(_13_), .Y(_13__bF_buf2) );
BUFX4 BUFX4_4 ( .A(_13_), .Y(_13__bF_buf1) );
BUFX4 BUFX4_5 ( .A(_13_), .Y(_13__bF_buf0) );
BUFX4 BUFX4_6 ( .A(_51_), .Y(_51__bF_buf5) );
BUFX4 BUFX4_7 ( .A(_51_), .Y(_51__bF_buf4) );
BUFX4 BUFX4_8 ( .A(_51_), .Y(_51__bF_buf3) );
BUFX4 BUFX4_9 ( .A(_51_), .Y(_51__bF_buf2) );
BUFX4 BUFX4_10 ( .A(_51_), .Y(_51__bF_buf1) );
BUFX4 BUFX4_11 ( .A(_51_), .Y(_51__bF_buf0) );
BUFX4 BUFX4_12 ( .A(_373_), .Y(_373__bF_buf3) );
BUFX4 BUFX4_13 ( .A(_373_), .Y(_373__bF_buf2) );
BUFX2 BUFX2_1 ( .A(_373_), .Y(_373__bF_buf1) );
BUFX4 BUFX4_14 ( .A(_373_), .Y(_373__bF_buf0) );
BUFX4 BUFX4_15 ( .A(_429_), .Y(_429__bF_buf7) );
BUFX4 BUFX4_16 ( .A(_429_), .Y(_429__bF_buf6) );
BUFX4 BUFX4_17 ( .A(_429_), .Y(_429__bF_buf5) );
BUFX4 BUFX4_18 ( .A(_429_), .Y(_429__bF_buf4) );
BUFX4 BUFX4_19 ( .A(_429_), .Y(_429__bF_buf3) );
BUFX4 BUFX4_20 ( .A(_429_), .Y(_429__bF_buf2) );
BUFX4 BUFX4_21 ( .A(_429_), .Y(_429__bF_buf1) );
BUFX4 BUFX4_22 ( .A(_429_), .Y(_429__bF_buf0) );
BUFX4 BUFX4_23 ( .A(CLK_I), .Y(CLK_I_bF_buf7) );
BUFX4 BUFX4_24 ( .A(CLK_I), .Y(CLK_I_bF_buf6) );
BUFX4 BUFX4_25 ( .A(CLK_I), .Y(CLK_I_bF_buf5) );
BUFX4 BUFX4_26 ( .A(CLK_I), .Y(CLK_I_bF_buf4) );
BUFX4 BUFX4_27 ( .A(CLK_I), .Y(CLK_I_bF_buf3) );
BUFX4 BUFX4_28 ( .A(CLK_I), .Y(CLK_I_bF_buf2) );
BUFX4 BUFX4_29 ( .A(CLK_I), .Y(CLK_I_bF_buf1) );
BUFX4 BUFX4_30 ( .A(CLK_I), .Y(CLK_I_bF_buf0) );
BUFX4 BUFX4_31 ( .A(status_1_), .Y(status_1_bF_buf3) );
BUFX4 BUFX4_32 ( .A(status_1_), .Y(status_1_bF_buf2) );
BUFX2 BUFX2_2 ( .A(status_1_), .Y(status_1_bF_buf1) );
BUFX2 BUFX2_3 ( .A(status_1_), .Y(status_1_bF_buf0) );
BUFX2 BUFX2_4 ( .A(status_0_), .Y(status_0_bF_buf3) );
BUFX2 BUFX2_5 ( .A(status_0_), .Y(status_0_bF_buf2) );
BUFX2 BUFX2_6 ( .A(status_0_), .Y(status_0_bF_buf1) );
BUFX2 BUFX2_7 ( .A(status_0_), .Y(status_0_bF_buf0) );
INVX2 INVX2_1 ( .A(reg_start), .Y(_12_) );
NOR2X1 NOR2X1_1 ( .A(reg_stop), .B(_12_), .Y(_13_) );
INVX4 INVX4_1 ( .A(dw08_cs), .Y(_15_) );
INVX4 INVX4_2 ( .A(reg_wr), .Y(_16_) );
OAI21X1 OAI21X1_1 ( .A(_15_), .B(_16_), .C(status_0_bF_buf1), .Y(_17_) );
INVX1 INVX1_1 ( .A(_17_), .Y(_18_) );
OAI21X1 OAI21X1_2 ( .A(status_1_bF_buf0), .B(_18_), .C(_13__bF_buf0), .Y(_19_) );
INVX1 INVX1_2 ( .A(internal_counter_11_), .Y(_20_) );
INVX2 INVX2_2 ( .A(internal_counter_8_), .Y(_21_) );
NOR2X1 NOR2X1_2 ( .A(internal_counter_10_), .B(internal_counter_9_), .Y(_22_) );
NAND3X1 NAND3X1_1 ( .A(_20_), .B(_21_), .C(_22_), .Y(_23_) );
INVX2 INVX2_3 ( .A(internal_counter_4_), .Y(_24_) );
INVX1 INVX1_3 ( .A(internal_counter_5_), .Y(_25_) );
NOR2X1 NOR2X1_3 ( .A(internal_counter_6_), .B(internal_counter_7_), .Y(_26_) );
NAND3X1 NAND3X1_2 ( .A(_24_), .B(_25_), .C(_26_), .Y(_27_) );
NOR2X1 NOR2X1_4 ( .A(_23_), .B(_27_), .Y(_28_) );
NOR2X1 NOR2X1_5 ( .A(internal_counter_0_), .B(internal_counter_1_), .Y(_29_) );
NOR2X1 NOR2X1_6 ( .A(internal_counter_2_), .B(internal_counter_3_), .Y(_30_) );
NAND2X1 NAND2X1_1 ( .A(_29_), .B(_30_), .Y(_32_) );
INVX1 INVX1_4 ( .A(internal_counter_14_), .Y(_33_) );
INVX2 INVX2_4 ( .A(internal_counter_15_), .Y(_34_) );
NOR2X1 NOR2X1_7 ( .A(internal_counter_12_), .B(internal_counter_13_), .Y(_35_) );
NAND3X1 NAND3X1_3 ( .A(_33_), .B(_34_), .C(_35_), .Y(_36_) );
NOR2X1 NOR2X1_8 ( .A(_32_), .B(_36_), .Y(_37_) );
NAND2X1 NAND2X1_2 ( .A(_37_), .B(_28_), .Y(_38_) );
INVX2 INVX2_5 ( .A(status_2_), .Y(_39_) );
INVX1 INVX1_5 ( .A(reg_stop), .Y(_40_) );
AND2X2 AND2X2_1 ( .A(_28_), .B(_37_), .Y(_41_) );
NOR2X1 NOR2X1_9 ( .A(_40_), .B(_41_), .Y(_42_) );
NOR2X1 NOR2X1_10 ( .A(_39_), .B(_42_), .Y(_43_) );
OAI21X1 OAI21X1_3 ( .A(reg_cont), .B(_38_), .C(_43_), .Y(_44_) );
NAND2X1 NAND2X1_3 ( .A(_19_), .B(_44_), .Y(_424__2_) );
INVX1 INVX1_6 ( .A(status_1_bF_buf1), .Y(_45_) );
NAND3X1 NAND3X1_4 ( .A(reg_stop), .B(status_2_), .C(_38_), .Y(_46_) );
OAI21X1 OAI21X1_4 ( .A(_45_), .B(_13__bF_buf1), .C(_46_), .Y(_424__1_) );
INVX1 INVX1_7 ( .A(reg_cont), .Y(_47_) );
NAND2X1 NAND2X1_4 ( .A(_47_), .B(_41_), .Y(_49_) );
INVX2 INVX2_6 ( .A(_13__bF_buf0), .Y(_50_) );
NOR2X1 NOR2X1_11 ( .A(_15_), .B(_16_), .Y(_51_) );
OAI21X1 OAI21X1_5 ( .A(_51__bF_buf1), .B(_50_), .C(status_0_bF_buf1), .Y(_52_) );
OAI21X1 OAI21X1_6 ( .A(_39_), .B(_49_), .C(_52_), .Y(_424__0_) );
INVX1 INVX1_8 ( .A(S_ADR_I[3]), .Y(_53_) );
NOR2X1 NOR2X1_12 ( .A(S_ADR_I[5]), .B(S_ADR_I[4]), .Y(_54_) );
NAND2X1 NAND2X1_5 ( .A(_53_), .B(_54_), .Y(_55_) );
NOR2X1 NOR2X1_13 ( .A(S_ADR_I[2]), .B(_55_), .Y(_0_) );
INVX1 INVX1_9 ( .A(S_ADR_I[2]), .Y(_56_) );
NOR2X1 NOR2X1_14 ( .A(_56_), .B(_55_), .Y(_1_) );
NAND2X1 NAND2X1_6 ( .A(S_ADR_I[3]), .B(_54_), .Y(_57_) );
NOR2X1 NOR2X1_15 ( .A(S_ADR_I[2]), .B(_57_), .Y(_2_) );
NOR2X1 NOR2X1_16 ( .A(_56_), .B(_57_), .Y(_3_) );
AND2X2 AND2X2_2 ( .A(S_STB_I), .B(S_CYC_I), .Y(_11_) );
NAND2X1 NAND2X1_7 ( .A(S_WE_I), .B(_11_), .Y(_58_) );
INVX1 INVX1_10 ( .A(_58_), .Y(_10_) );
NAND2X1 NAND2X1_8 ( .A(reg_run), .B(_41_), .Y(_59_) );
NOR2X1 NOR2X1_17 ( .A(_428_), .B(_59_), .Y(_423_) );
NAND2X1 NAND2X1_9 ( .A(latch_s_data_0_), .B(_51__bF_buf5), .Y(_61_) );
INVX1 INVX1_11 ( .A(_61_), .Y(_62_) );
INVX2 INVX2_7 ( .A(internal_counter_0_), .Y(_63_) );
NOR2X1 NOR2X1_18 ( .A(reg_08_data_10_), .B(reg_08_data_11_), .Y(_64_) );
NOR2X1 NOR2X1_19 ( .A(reg_08_data_8_), .B(reg_08_data_9_), .Y(_65_) );
NAND2X1 NAND2X1_10 ( .A(_64_), .B(_65_), .Y(_66_) );
NOR2X1 NOR2X1_20 ( .A(reg_08_data_6_), .B(reg_08_data_7_), .Y(_67_) );
NOR2X1 NOR2X1_21 ( .A(reg_08_data_4_), .B(reg_08_data_5_), .Y(_68_) );
NAND2X1 NAND2X1_11 ( .A(_67_), .B(_68_), .Y(_69_) );
NOR2X1 NOR2X1_22 ( .A(_66_), .B(_69_), .Y(_70_) );
NOR2X1 NOR2X1_23 ( .A(reg_08_data_0_), .B(reg_08_data_1_), .Y(_71_) );
NOR2X1 NOR2X1_24 ( .A(reg_08_data_2_), .B(reg_08_data_3_), .Y(_72_) );
NAND2X1 NAND2X1_12 ( .A(_71_), .B(_72_), .Y(_73_) );
INVX1 INVX1_12 ( .A(reg_08_data_14_), .Y(_74_) );
INVX1 INVX1_13 ( .A(reg_08_data_15_), .Y(_75_) );
NOR2X1 NOR2X1_25 ( .A(reg_08_data_12_), .B(reg_08_data_13_), .Y(_76_) );
NAND3X1 NAND3X1_5 ( .A(_74_), .B(_75_), .C(_76_), .Y(_77_) );
NOR2X1 NOR2X1_26 ( .A(_73_), .B(_77_), .Y(_78_) );
NAND2X1 NAND2X1_13 ( .A(_70_), .B(_78_), .Y(_79_) );
NAND2X1 NAND2X1_14 ( .A(_13__bF_buf4), .B(_79_), .Y(_80_) );
INVX1 INVX1_14 ( .A(reg_08_data_0_), .Y(_82_) );
INVX4 INVX4_3 ( .A(_51__bF_buf3), .Y(_83_) );
OAI21X1 OAI21X1_7 ( .A(_82_), .B(_50_), .C(_83_), .Y(_84_) );
AOI21X1 AOI21X1_1 ( .A(_80_), .B(_63_), .C(_84_), .Y(_85_) );
OAI21X1 OAI21X1_8 ( .A(_62_), .B(_85_), .C(status_0_bF_buf3), .Y(_86_) );
NAND2X1 NAND2X1_15 ( .A(_63_), .B(_38_), .Y(_87_) );
NAND2X1 NAND2X1_16 ( .A(reg_08_data_0_), .B(_41_), .Y(_88_) );
AOI21X1 AOI21X1_2 ( .A(_88_), .B(_87_), .C(_51__bF_buf5), .Y(_89_) );
OAI21X1 OAI21X1_9 ( .A(_62_), .B(_89_), .C(_43_), .Y(_90_) );
INVX4 INVX4_4 ( .A(_46_), .Y(_91_) );
OAI21X1 OAI21X1_10 ( .A(reg_stop), .B(_12_), .C(_51__bF_buf1), .Y(_92_) );
INVX4 INVX4_5 ( .A(_92_), .Y(_93_) );
OAI22X1 OAI22X1_1 ( .A(_13__bF_buf2), .B(_61_), .C(_63_), .D(_93_), .Y(_94_) );
AOI22X1 AOI22X1_1 ( .A(status_1_bF_buf2), .B(_94_), .C(internal_counter_0_), .D(_91_), .Y(_95_) );
NAND3X1 NAND3X1_6 ( .A(_86_), .B(_95_), .C(_90_), .Y(_14_) );
NAND2X1 NAND2X1_17 ( .A(latch_s_data_1_), .B(_51__bF_buf5), .Y(_96_) );
INVX1 INVX1_15 ( .A(_96_), .Y(_97_) );
INVX2 INVX2_8 ( .A(internal_counter_1_), .Y(_98_) );
INVX1 INVX1_16 ( .A(reg_08_data_1_), .Y(_100_) );
NOR2X1 NOR2X1_27 ( .A(_82_), .B(_100_), .Y(_101_) );
OAI21X1 OAI21X1_11 ( .A(reg_08_data_0_), .B(reg_08_data_1_), .C(_13__bF_buf2), .Y(_102_) );
OAI21X1 OAI21X1_12 ( .A(_101_), .B(_102_), .C(_83_), .Y(_103_) );
AOI21X1 AOI21X1_3 ( .A(_80_), .B(_98_), .C(_103_), .Y(_104_) );
OAI21X1 OAI21X1_13 ( .A(_97_), .B(_104_), .C(status_0_bF_buf3), .Y(_105_) );
NOR2X1 NOR2X1_28 ( .A(_63_), .B(_98_), .Y(_106_) );
OAI21X1 OAI21X1_14 ( .A(_29_), .B(_106_), .C(_38_), .Y(_107_) );
NAND2X1 NAND2X1_18 ( .A(reg_08_data_1_), .B(_41_), .Y(_108_) );
AOI21X1 AOI21X1_4 ( .A(_108_), .B(_107_), .C(_51__bF_buf3), .Y(_109_) );
OAI21X1 OAI21X1_15 ( .A(_97_), .B(_109_), .C(_43_), .Y(_110_) );
OAI22X1 OAI22X1_2 ( .A(_13__bF_buf2), .B(_96_), .C(_98_), .D(_93_), .Y(_111_) );
AOI22X1 AOI22X1_2 ( .A(status_1_bF_buf2), .B(_111_), .C(internal_counter_1_), .D(_91_), .Y(_112_) );
NAND3X1 NAND3X1_7 ( .A(_105_), .B(_112_), .C(_110_), .Y(_31_) );
NAND2X1 NAND2X1_19 ( .A(latch_s_data_2_), .B(_51__bF_buf3), .Y(_113_) );
INVX1 INVX1_17 ( .A(_113_), .Y(_114_) );
INVX1 INVX1_18 ( .A(internal_counter_2_), .Y(_115_) );
OAI21X1 OAI21X1_16 ( .A(reg_08_data_0_), .B(reg_08_data_1_), .C(reg_08_data_2_), .Y(_116_) );
INVX1 INVX1_19 ( .A(_116_), .Y(_117_) );
INVX1 INVX1_20 ( .A(_71_), .Y(_118_) );
OAI21X1 OAI21X1_17 ( .A(reg_08_data_2_), .B(_118_), .C(_13__bF_buf2), .Y(_119_) );
OAI21X1 OAI21X1_18 ( .A(_117_), .B(_119_), .C(_83_), .Y(_121_) );
AOI21X1 AOI21X1_5 ( .A(_80_), .B(_115_), .C(_121_), .Y(_122_) );
OAI21X1 OAI21X1_19 ( .A(_114_), .B(_122_), .C(status_0_bF_buf3), .Y(_123_) );
NAND2X1 NAND2X1_20 ( .A(_115_), .B(_29_), .Y(_124_) );
OAI21X1 OAI21X1_20 ( .A(internal_counter_0_), .B(internal_counter_1_), .C(internal_counter_2_), .Y(_125_) );
NAND2X1 NAND2X1_21 ( .A(_125_), .B(_124_), .Y(_126_) );
OAI21X1 OAI21X1_21 ( .A(reg_08_data_2_), .B(_38_), .C(_126_), .Y(_127_) );
OAI21X1 OAI21X1_22 ( .A(_51__bF_buf3), .B(_127_), .C(_113_), .Y(_128_) );
NAND2X1 NAND2X1_22 ( .A(_128_), .B(_43_), .Y(_129_) );
OAI22X1 OAI22X1_3 ( .A(_13__bF_buf4), .B(_113_), .C(_115_), .D(_93_), .Y(_130_) );
AOI22X1 AOI22X1_3 ( .A(status_1_bF_buf2), .B(_130_), .C(internal_counter_2_), .D(_91_), .Y(_131_) );
NAND3X1 NAND3X1_8 ( .A(_131_), .B(_123_), .C(_129_), .Y(_48_) );
NAND2X1 NAND2X1_23 ( .A(latch_s_data_3_), .B(_51__bF_buf5), .Y(_132_) );
INVX1 INVX1_21 ( .A(_132_), .Y(_133_) );
INVX2 INVX2_9 ( .A(internal_counter_3_), .Y(_134_) );
INVX1 INVX1_22 ( .A(reg_08_data_2_), .Y(_135_) );
INVX1 INVX1_23 ( .A(reg_08_data_3_), .Y(_136_) );
AOI21X1 AOI21X1_6 ( .A(_71_), .B(_135_), .C(_136_), .Y(_137_) );
NAND2X1 NAND2X1_24 ( .A(_13__bF_buf4), .B(_73_), .Y(_139_) );
OAI21X1 OAI21X1_23 ( .A(_137_), .B(_139_), .C(_83_), .Y(_140_) );
AOI21X1 AOI21X1_7 ( .A(_80_), .B(_134_), .C(_140_), .Y(_141_) );
OAI21X1 OAI21X1_24 ( .A(_133_), .B(_141_), .C(status_0_bF_buf3), .Y(_142_) );
XNOR2X1 XNOR2X1_1 ( .A(_124_), .B(_134_), .Y(_143_) );
OAI21X1 OAI21X1_25 ( .A(reg_08_data_3_), .B(_38_), .C(_83_), .Y(_144_) );
OAI21X1 OAI21X1_26 ( .A(_143_), .B(_144_), .C(_132_), .Y(_145_) );
NAND2X1 NAND2X1_25 ( .A(_145_), .B(_43_), .Y(_146_) );
OAI22X1 OAI22X1_4 ( .A(_13__bF_buf2), .B(_132_), .C(_134_), .D(_93_), .Y(_147_) );
AOI22X1 AOI22X1_4 ( .A(status_1_bF_buf2), .B(_147_), .C(internal_counter_3_), .D(_91_), .Y(_148_) );
NAND3X1 NAND3X1_9 ( .A(_148_), .B(_142_), .C(_146_), .Y(_60_) );
NAND2X1 NAND2X1_26 ( .A(latch_s_data_4_), .B(_51__bF_buf4), .Y(_149_) );
INVX1 INVX1_24 ( .A(_149_), .Y(_150_) );
INVX1 INVX1_25 ( .A(reg_08_data_4_), .Y(_151_) );
AND2X2 AND2X2_3 ( .A(_71_), .B(_72_), .Y(_152_) );
NOR2X1 NOR2X1_29 ( .A(_151_), .B(_152_), .Y(_153_) );
OAI21X1 OAI21X1_27 ( .A(reg_08_data_4_), .B(_73_), .C(_13__bF_buf4), .Y(_154_) );
OAI21X1 OAI21X1_28 ( .A(_154_), .B(_153_), .C(_83_), .Y(_155_) );
AOI21X1 AOI21X1_8 ( .A(_80_), .B(_24_), .C(_155_), .Y(_156_) );
OAI21X1 OAI21X1_29 ( .A(_150_), .B(_156_), .C(status_0_bF_buf0), .Y(_157_) );
NOR2X1 NOR2X1_30 ( .A(_24_), .B(_93_), .Y(_158_) );
NOR2X1 NOR2X1_31 ( .A(_13__bF_buf4), .B(_149_), .Y(_159_) );
OAI21X1 OAI21X1_30 ( .A(_159_), .B(_158_), .C(status_1_bF_buf1), .Y(_160_) );
NAND3X1 NAND3X1_10 ( .A(_24_), .B(_29_), .C(_30_), .Y(_162_) );
OAI21X1 OAI21X1_31 ( .A(internal_counter_3_), .B(_124_), .C(internal_counter_4_), .Y(_163_) );
OAI21X1 OAI21X1_32 ( .A(reg_08_data_4_), .B(_38_), .C(_83_), .Y(_164_) );
AOI21X1 AOI21X1_9 ( .A(_162_), .B(_163_), .C(_164_), .Y(_165_) );
OAI21X1 OAI21X1_33 ( .A(_40_), .B(_41_), .C(_149_), .Y(_166_) );
AOI21X1 AOI21X1_10 ( .A(_42_), .B(_24_), .C(_39_), .Y(_167_) );
OAI21X1 OAI21X1_34 ( .A(_165_), .B(_166_), .C(_167_), .Y(_168_) );
NAND3X1 NAND3X1_11 ( .A(_157_), .B(_160_), .C(_168_), .Y(_81_) );
AOI21X1 AOI21X1_11 ( .A(_78_), .B(_70_), .C(_50_), .Y(_169_) );
OAI21X1 OAI21X1_35 ( .A(reg_08_data_4_), .B(_73_), .C(reg_08_data_5_), .Y(_170_) );
NAND3X1 NAND3X1_12 ( .A(_68_), .B(_71_), .C(_72_), .Y(_171_) );
INVX1 INVX1_26 ( .A(_171_), .Y(_172_) );
NOR2X1 NOR2X1_32 ( .A(_50_), .B(_172_), .Y(_173_) );
AOI21X1 AOI21X1_12 ( .A(_173_), .B(_170_), .C(_17_), .Y(_174_) );
OAI21X1 OAI21X1_36 ( .A(internal_counter_5_), .B(_169_), .C(_174_), .Y(_175_) );
NAND2X1 NAND2X1_27 ( .A(latch_s_data_5_), .B(_51__bF_buf1), .Y(_176_) );
NOR2X1 NOR2X1_33 ( .A(internal_counter_5_), .B(_162_), .Y(_177_) );
AND2X2 AND2X2_4 ( .A(_162_), .B(internal_counter_5_), .Y(_178_) );
OAI22X1 OAI22X1_5 ( .A(_177_), .B(_178_), .C(reg_08_data_5_), .D(_38_), .Y(_180_) );
OAI21X1 OAI21X1_37 ( .A(_51__bF_buf2), .B(_180_), .C(_176_), .Y(_181_) );
NAND2X1 NAND2X1_28 ( .A(_181_), .B(_43_), .Y(_182_) );
NAND3X1 NAND3X1_13 ( .A(internal_counter_5_), .B(status_1_bF_buf1), .C(_92_), .Y(_183_) );
OAI21X1 OAI21X1_38 ( .A(reg_stop), .B(_12_), .C(status_1_bF_buf0), .Y(_184_) );
INVX1 INVX1_27 ( .A(_184_), .Y(_185_) );
NOR2X1 NOR2X1_34 ( .A(status_0_bF_buf0), .B(_185_), .Y(_186_) );
OAI21X1 OAI21X1_39 ( .A(_176_), .B(_186_), .C(_183_), .Y(_187_) );
AOI21X1 AOI21X1_13 ( .A(_91_), .B(internal_counter_5_), .C(_187_), .Y(_188_) );
NAND3X1 NAND3X1_14 ( .A(_175_), .B(_188_), .C(_182_), .Y(_99_) );
NAND2X1 NAND2X1_29 ( .A(latch_s_data_6_), .B(_51__bF_buf4), .Y(_189_) );
INVX1 INVX1_28 ( .A(_189_), .Y(_190_) );
INVX1 INVX1_29 ( .A(internal_counter_6_), .Y(_191_) );
NOR2X1 NOR2X1_35 ( .A(reg_08_data_6_), .B(_171_), .Y(_192_) );
INVX1 INVX1_30 ( .A(reg_08_data_6_), .Y(_193_) );
OAI21X1 OAI21X1_40 ( .A(_193_), .B(_172_), .C(_13__bF_buf1), .Y(_194_) );
OAI21X1 OAI21X1_41 ( .A(_192_), .B(_194_), .C(_83_), .Y(_195_) );
AOI21X1 AOI21X1_14 ( .A(_191_), .B(_80_), .C(_195_), .Y(_196_) );
OAI21X1 OAI21X1_42 ( .A(_190_), .B(_196_), .C(status_0_bF_buf0), .Y(_197_) );
NAND2X1 NAND2X1_30 ( .A(_191_), .B(_25_), .Y(_198_) );
OAI21X1 OAI21X1_43 ( .A(internal_counter_5_), .B(_162_), .C(internal_counter_6_), .Y(_199_) );
OAI21X1 OAI21X1_44 ( .A(_162_), .B(_198_), .C(_199_), .Y(_200_) );
OAI21X1 OAI21X1_45 ( .A(reg_08_data_6_), .B(_38_), .C(_200_), .Y(_201_) );
OAI21X1 OAI21X1_46 ( .A(_51__bF_buf4), .B(_201_), .C(_189_), .Y(_202_) );
NAND2X1 NAND2X1_31 ( .A(_202_), .B(_43_), .Y(_203_) );
OAI21X1 OAI21X1_47 ( .A(_45_), .B(_93_), .C(_46_), .Y(_205_) );
AOI22X1 AOI22X1_5 ( .A(_185_), .B(_190_), .C(internal_counter_6_), .D(_205_), .Y(_206_) );
NAND3X1 NAND3X1_15 ( .A(_206_), .B(_203_), .C(_197_), .Y(_120_) );
NAND2X1 NAND2X1_32 ( .A(latch_s_data_7_), .B(_51__bF_buf4), .Y(_207_) );
NOR2X1 NOR2X1_36 ( .A(_73_), .B(_69_), .Y(_208_) );
INVX1 INVX1_31 ( .A(reg_08_data_7_), .Y(_209_) );
OAI21X1 OAI21X1_48 ( .A(_209_), .B(_192_), .C(_13__bF_buf1), .Y(_210_) );
OAI22X1 OAI22X1_6 ( .A(internal_counter_7_), .B(_169_), .C(_208_), .D(_210_), .Y(_211_) );
OAI21X1 OAI21X1_49 ( .A(_51__bF_buf2), .B(_211_), .C(_207_), .Y(_212_) );
NAND2X1 NAND2X1_33 ( .A(status_0_bF_buf0), .B(_212_), .Y(_213_) );
INVX1 INVX1_32 ( .A(_207_), .Y(_214_) );
AND2X2 AND2X2_5 ( .A(internal_counter_7_), .B(status_1_bF_buf1), .Y(_215_) );
AOI22X1 AOI22X1_6 ( .A(_92_), .B(_215_), .C(_185_), .D(_214_), .Y(_216_) );
NAND2X1 NAND2X1_34 ( .A(_25_), .B(_26_), .Y(_217_) );
OAI21X1 OAI21X1_50 ( .A(_198_), .B(_162_), .C(internal_counter_7_), .Y(_218_) );
OAI21X1 OAI21X1_51 ( .A(_162_), .B(_217_), .C(_218_), .Y(_219_) );
OAI21X1 OAI21X1_52 ( .A(reg_08_data_7_), .B(_38_), .C(_219_), .Y(_220_) );
OAI21X1 OAI21X1_53 ( .A(_51__bF_buf2), .B(_220_), .C(_207_), .Y(_221_) );
AOI22X1 AOI22X1_7 ( .A(internal_counter_7_), .B(_91_), .C(_221_), .D(_43_), .Y(_223_) );
NAND3X1 NAND3X1_16 ( .A(_216_), .B(_223_), .C(_213_), .Y(_138_) );
NAND2X1 NAND2X1_35 ( .A(latch_s_data_8_), .B(_51__bF_buf2), .Y(_224_) );
INVX2 INVX2_10 ( .A(reg_08_data_8_), .Y(_225_) );
AND2X2 AND2X2_6 ( .A(_208_), .B(_225_), .Y(_226_) );
OAI21X1 OAI21X1_54 ( .A(_225_), .B(_208_), .C(_13__bF_buf1), .Y(_227_) );
OAI22X1 OAI22X1_7 ( .A(_226_), .B(_227_), .C(internal_counter_8_), .D(_169_), .Y(_228_) );
OAI21X1 OAI21X1_55 ( .A(_51__bF_buf0), .B(_228_), .C(_224_), .Y(_229_) );
NAND2X1 NAND2X1_36 ( .A(status_0_bF_buf2), .B(_229_), .Y(_230_) );
OAI22X1 OAI22X1_8 ( .A(_13__bF_buf1), .B(_224_), .C(_21_), .D(_93_), .Y(_231_) );
NAND2X1 NAND2X1_37 ( .A(status_1_bF_buf3), .B(_231_), .Y(_232_) );
OAI21X1 OAI21X1_56 ( .A(_217_), .B(_162_), .C(internal_counter_8_), .Y(_233_) );
NOR2X1 NOR2X1_37 ( .A(_217_), .B(_162_), .Y(_234_) );
NAND2X1 NAND2X1_38 ( .A(_21_), .B(_234_), .Y(_235_) );
AND2X2 AND2X2_7 ( .A(_235_), .B(_233_), .Y(_236_) );
OAI21X1 OAI21X1_57 ( .A(reg_08_data_8_), .B(_38_), .C(_83_), .Y(_237_) );
OAI21X1 OAI21X1_58 ( .A(_236_), .B(_237_), .C(_224_), .Y(_238_) );
AOI22X1 AOI22X1_8 ( .A(internal_counter_8_), .B(_91_), .C(_238_), .D(_43_), .Y(_239_) );
NAND3X1 NAND3X1_17 ( .A(_232_), .B(_230_), .C(_239_), .Y(_161_) );
NAND2X1 NAND2X1_39 ( .A(latch_s_data_9_), .B(_51__bF_buf0), .Y(_240_) );
INVX1 INVX1_33 ( .A(reg_08_data_9_), .Y(_241_) );
AOI21X1 AOI21X1_15 ( .A(_208_), .B(_225_), .C(_241_), .Y(_242_) );
AND2X2 AND2X2_8 ( .A(_67_), .B(_68_), .Y(_244_) );
NAND3X1 NAND3X1_18 ( .A(_65_), .B(_244_), .C(_152_), .Y(_245_) );
NAND2X1 NAND2X1_40 ( .A(_13__bF_buf3), .B(_245_), .Y(_246_) );
OAI22X1 OAI22X1_9 ( .A(_246_), .B(_242_), .C(internal_counter_9_), .D(_169_), .Y(_247_) );
OAI21X1 OAI21X1_59 ( .A(_51__bF_buf0), .B(_247_), .C(_240_), .Y(_248_) );
NAND2X1 NAND2X1_41 ( .A(status_0_bF_buf2), .B(_248_), .Y(_249_) );
INVX1 INVX1_34 ( .A(_240_), .Y(_250_) );
INVX1 INVX1_35 ( .A(internal_counter_9_), .Y(_251_) );
NAND3X1 NAND3X1_19 ( .A(_21_), .B(_251_), .C(_234_), .Y(_252_) );
INVX1 INVX1_36 ( .A(_234_), .Y(_253_) );
OAI21X1 OAI21X1_60 ( .A(internal_counter_8_), .B(_253_), .C(internal_counter_9_), .Y(_254_) );
OAI21X1 OAI21X1_61 ( .A(reg_08_data_9_), .B(_38_), .C(_83_), .Y(_255_) );
AOI21X1 AOI21X1_16 ( .A(_254_), .B(_252_), .C(_255_), .Y(_256_) );
OAI21X1 OAI21X1_62 ( .A(_250_), .B(_256_), .C(_43_), .Y(_257_) );
OAI22X1 OAI22X1_10 ( .A(_13__bF_buf3), .B(_240_), .C(_251_), .D(_93_), .Y(_258_) );
AOI22X1 AOI22X1_9 ( .A(status_1_bF_buf3), .B(_258_), .C(internal_counter_9_), .D(_91_), .Y(_259_) );
NAND3X1 NAND3X1_20 ( .A(_259_), .B(_257_), .C(_249_), .Y(_179_) );
NAND2X1 NAND2X1_42 ( .A(latch_s_data_10_), .B(_51__bF_buf0), .Y(_260_) );
INVX1 INVX1_37 ( .A(reg_08_data_10_), .Y(_262_) );
AOI21X1 AOI21X1_17 ( .A(_208_), .B(_65_), .C(_262_), .Y(_263_) );
OAI21X1 OAI21X1_63 ( .A(reg_08_data_10_), .B(_245_), .C(_13__bF_buf3), .Y(_264_) );
OAI22X1 OAI22X1_11 ( .A(internal_counter_10_), .B(_169_), .C(_263_), .D(_264_), .Y(_265_) );
OAI21X1 OAI21X1_64 ( .A(_51__bF_buf0), .B(_265_), .C(_260_), .Y(_266_) );
NAND2X1 NAND2X1_43 ( .A(status_0_bF_buf2), .B(_266_), .Y(_267_) );
INVX1 INVX1_38 ( .A(_260_), .Y(_268_) );
OAI21X1 OAI21X1_65 ( .A(internal_counter_9_), .B(_235_), .C(internal_counter_10_), .Y(_269_) );
NAND3X1 NAND3X1_21 ( .A(_21_), .B(_22_), .C(_234_), .Y(_270_) );
OAI21X1 OAI21X1_66 ( .A(reg_08_data_10_), .B(_38_), .C(_83_), .Y(_271_) );
AOI21X1 AOI21X1_18 ( .A(_269_), .B(_270_), .C(_271_), .Y(_272_) );
OAI21X1 OAI21X1_67 ( .A(_268_), .B(_272_), .C(_43_), .Y(_273_) );
NAND3X1 NAND3X1_22 ( .A(internal_counter_10_), .B(status_1_bF_buf3), .C(_92_), .Y(_274_) );
OAI21X1 OAI21X1_68 ( .A(_184_), .B(_260_), .C(_274_), .Y(_275_) );
AOI21X1 AOI21X1_19 ( .A(_91_), .B(internal_counter_10_), .C(_275_), .Y(_276_) );
NAND3X1 NAND3X1_23 ( .A(_276_), .B(_273_), .C(_267_), .Y(_204_) );
OAI21X1 OAI21X1_69 ( .A(internal_counter_10_), .B(_252_), .C(internal_counter_11_), .Y(_277_) );
NOR3X1 NOR3X1_1 ( .A(_217_), .B(_23_), .C(_162_), .Y(_278_) );
AOI22X1 AOI22X1_10 ( .A(_36_), .B(_278_), .C(reg_08_data_11_), .D(_41_), .Y(_279_) );
NAND2X1 NAND2X1_44 ( .A(_277_), .B(_279_), .Y(_280_) );
NAND2X1 NAND2X1_45 ( .A(_20_), .B(_80_), .Y(_281_) );
INVX1 INVX1_39 ( .A(status_0_bF_buf1), .Y(_282_) );
OAI21X1 OAI21X1_70 ( .A(reg_08_data_10_), .B(_245_), .C(reg_08_data_11_), .Y(_283_) );
NOR3X1 NOR3X1_2 ( .A(_73_), .B(_66_), .C(_69_), .Y(_284_) );
NOR2X1 NOR2X1_38 ( .A(_50_), .B(_284_), .Y(_285_) );
AOI21X1 AOI21X1_20 ( .A(_285_), .B(_283_), .C(_282_), .Y(_286_) );
AOI22X1 AOI22X1_11 ( .A(_281_), .B(_286_), .C(_280_), .D(_43_), .Y(_287_) );
NAND2X1 NAND2X1_46 ( .A(latch_s_data_11_), .B(_51__bF_buf4), .Y(_288_) );
INVX1 INVX1_40 ( .A(_288_), .Y(_289_) );
OAI21X1 OAI21X1_71 ( .A(_39_), .B(_42_), .C(_186_), .Y(_290_) );
AOI22X1 AOI22X1_12 ( .A(internal_counter_11_), .B(_205_), .C(_289_), .D(_290_), .Y(_291_) );
OAI21X1 OAI21X1_72 ( .A(_51__bF_buf2), .B(_287_), .C(_291_), .Y(_222_) );
INVX1 INVX1_41 ( .A(reg_08_data_12_), .Y(_292_) );
NOR2X1 NOR2X1_39 ( .A(_292_), .B(_284_), .Y(_293_) );
AND2X2 AND2X2_9 ( .A(_64_), .B(_65_), .Y(_294_) );
NAND3X1 NAND3X1_24 ( .A(_294_), .B(_244_), .C(_152_), .Y(_295_) );
OAI21X1 OAI21X1_73 ( .A(reg_08_data_12_), .B(_295_), .C(_13__bF_buf0), .Y(_296_) );
OAI22X1 OAI22X1_12 ( .A(internal_counter_12_), .B(_169_), .C(_296_), .D(_293_), .Y(_297_) );
OAI21X1 OAI21X1_74 ( .A(_15_), .B(_16_), .C(_297_), .Y(_298_) );
OR2X2 OR2X2_1 ( .A(_83_), .B(latch_s_data_12_), .Y(_299_) );
NAND3X1 NAND3X1_25 ( .A(status_0_bF_buf1), .B(_299_), .C(_298_), .Y(_300_) );
NAND2X1 NAND2X1_47 ( .A(latch_s_data_12_), .B(_51__bF_buf1), .Y(_301_) );
INVX1 INVX1_42 ( .A(_301_), .Y(_302_) );
OAI21X1 OAI21X1_75 ( .A(_23_), .B(_253_), .C(internal_counter_12_), .Y(_303_) );
INVX2 INVX2_11 ( .A(internal_counter_12_), .Y(_304_) );
NAND2X1 NAND2X1_48 ( .A(_304_), .B(_278_), .Y(_305_) );
OAI21X1 OAI21X1_76 ( .A(reg_08_data_12_), .B(_38_), .C(_83_), .Y(_306_) );
AOI21X1 AOI21X1_21 ( .A(_303_), .B(_305_), .C(_306_), .Y(_307_) );
OAI21X1 OAI21X1_77 ( .A(_302_), .B(_307_), .C(_43_), .Y(_308_) );
OAI22X1 OAI22X1_13 ( .A(_13__bF_buf3), .B(_301_), .C(_304_), .D(_93_), .Y(_309_) );
AOI22X1 AOI22X1_13 ( .A(status_1_bF_buf3), .B(_309_), .C(internal_counter_12_), .D(_91_), .Y(_310_) );
NAND3X1 NAND3X1_26 ( .A(_308_), .B(_310_), .C(_300_), .Y(_243_) );
NOR2X1 NOR2X1_40 ( .A(internal_counter_13_), .B(_169_), .Y(_311_) );
NAND3X1 NAND3X1_27 ( .A(_292_), .B(_294_), .C(_208_), .Y(_312_) );
INVX1 INVX1_43 ( .A(_76_), .Y(_313_) );
OAI21X1 OAI21X1_78 ( .A(_313_), .B(_295_), .C(_13__bF_buf0), .Y(_314_) );
AOI21X1 AOI21X1_22 ( .A(reg_08_data_13_), .B(_312_), .C(_314_), .Y(_315_) );
OAI21X1 OAI21X1_79 ( .A(_311_), .B(_315_), .C(_83_), .Y(_316_) );
OR2X2 OR2X2_2 ( .A(_83_), .B(latch_s_data_13_), .Y(_317_) );
NAND3X1 NAND3X1_28 ( .A(status_0_bF_buf2), .B(_317_), .C(_316_), .Y(_318_) );
NAND2X1 NAND2X1_49 ( .A(latch_s_data_13_), .B(_51__bF_buf0), .Y(_319_) );
INVX1 INVX1_44 ( .A(_319_), .Y(_320_) );
OAI21X1 OAI21X1_80 ( .A(_15_), .B(_16_), .C(_38_), .Y(_321_) );
INVX1 INVX1_45 ( .A(internal_counter_13_), .Y(_322_) );
NAND3X1 NAND3X1_29 ( .A(_304_), .B(_322_), .C(_278_), .Y(_323_) );
NAND2X1 NAND2X1_50 ( .A(internal_counter_13_), .B(_305_), .Y(_324_) );
OAI21X1 OAI21X1_81 ( .A(_15_), .B(_16_), .C(reg_08_data_13_), .Y(_325_) );
AOI22X1 AOI22X1_14 ( .A(_321_), .B(_325_), .C(_323_), .D(_324_), .Y(_326_) );
OAI21X1 OAI21X1_82 ( .A(_320_), .B(_326_), .C(_43_), .Y(_327_) );
OAI22X1 OAI22X1_14 ( .A(_13__bF_buf3), .B(_319_), .C(_322_), .D(_93_), .Y(_328_) );
AOI22X1 AOI22X1_15 ( .A(status_1_bF_buf3), .B(_328_), .C(internal_counter_13_), .D(_91_), .Y(_329_) );
NAND3X1 NAND3X1_30 ( .A(_327_), .B(_329_), .C(_318_), .Y(_261_) );
NAND2X1 NAND2X1_51 ( .A(latch_s_data_14_), .B(_51__bF_buf1), .Y(_330_) );
INVX1 INVX1_46 ( .A(_330_), .Y(_331_) );
NAND2X1 NAND2X1_52 ( .A(internal_counter_14_), .B(_323_), .Y(_332_) );
NOR2X1 NOR2X1_41 ( .A(internal_counter_13_), .B(internal_counter_14_), .Y(_333_) );
NAND3X1 NAND3X1_31 ( .A(_304_), .B(_333_), .C(_278_), .Y(_334_) );
OAI21X1 OAI21X1_83 ( .A(_15_), .B(_16_), .C(reg_08_data_14_), .Y(_335_) );
AOI22X1 AOI22X1_16 ( .A(_321_), .B(_335_), .C(_334_), .D(_332_), .Y(_336_) );
OAI21X1 OAI21X1_84 ( .A(_331_), .B(_336_), .C(_43_), .Y(_337_) );
NAND2X1 NAND2X1_53 ( .A(_33_), .B(_80_), .Y(_338_) );
NAND3X1 NAND3X1_32 ( .A(_74_), .B(_76_), .C(_284_), .Y(_339_) );
OAI21X1 OAI21X1_85 ( .A(_313_), .B(_295_), .C(reg_08_data_14_), .Y(_340_) );
NAND3X1 NAND3X1_33 ( .A(_13__bF_buf0), .B(_339_), .C(_340_), .Y(_341_) );
NAND3X1 NAND3X1_34 ( .A(_18_), .B(_338_), .C(_341_), .Y(_342_) );
NAND3X1 NAND3X1_35 ( .A(internal_counter_14_), .B(status_1_bF_buf0), .C(_92_), .Y(_343_) );
OAI21X1 OAI21X1_86 ( .A(_330_), .B(_186_), .C(_343_), .Y(_344_) );
AOI21X1 AOI21X1_23 ( .A(_91_), .B(internal_counter_14_), .C(_344_), .Y(_345_) );
NAND3X1 NAND3X1_36 ( .A(_342_), .B(_345_), .C(_337_), .Y(_4__14_) );
NOR2X1 NOR2X1_42 ( .A(internal_counter_15_), .B(_169_), .Y(_346_) );
NOR2X1 NOR2X1_43 ( .A(_75_), .B(_51__bF_buf5), .Y(_347_) );
NAND2X1 NAND2X1_54 ( .A(_347_), .B(_339_), .Y(_348_) );
NOR2X1 NOR2X1_44 ( .A(_34_), .B(_51__bF_buf5), .Y(_349_) );
AOI22X1 AOI22X1_17 ( .A(latch_s_data_15_), .B(_51__bF_buf3), .C(_349_), .D(_80_), .Y(_350_) );
OAI21X1 OAI21X1_87 ( .A(_346_), .B(_348_), .C(_350_), .Y(_351_) );
NAND2X1 NAND2X1_55 ( .A(status_0_bF_buf3), .B(_351_), .Y(_352_) );
NOR2X1 NOR2X1_45 ( .A(_34_), .B(_93_), .Y(_353_) );
NAND2X1 NAND2X1_56 ( .A(latch_s_data_15_), .B(_51__bF_buf3), .Y(_354_) );
NOR2X1 NOR2X1_46 ( .A(_13__bF_buf4), .B(_354_), .Y(_355_) );
OAI21X1 OAI21X1_88 ( .A(_355_), .B(_353_), .C(status_1_bF_buf2), .Y(_356_) );
AND2X2 AND2X2_10 ( .A(_334_), .B(_349_), .Y(_357_) );
NAND2X1 NAND2X1_57 ( .A(reg_stop), .B(_38_), .Y(_358_) );
NAND2X1 NAND2X1_58 ( .A(_347_), .B(_41_), .Y(_359_) );
NAND3X1 NAND3X1_37 ( .A(_358_), .B(_354_), .C(_359_), .Y(_360_) );
AOI21X1 AOI21X1_24 ( .A(_42_), .B(_34_), .C(_39_), .Y(_361_) );
OAI21X1 OAI21X1_89 ( .A(_357_), .B(_360_), .C(_361_), .Y(_362_) );
NAND3X1 NAND3X1_38 ( .A(_356_), .B(_362_), .C(_352_), .Y(_4__15_) );
INVX1 INVX1_47 ( .A(_427_), .Y(_364_) );
INVX1 INVX1_48 ( .A(S_STB_I), .Y(_366_) );
NOR2X1 NOR2X1_47 ( .A(S_WE_I), .B(_366_), .Y(_368_) );
NAND2X1 NAND2X1_59 ( .A(dw00_cs), .B(_368_), .Y(_370_) );
INVX1 INVX1_49 ( .A(_368_), .Y(_372_) );
NOR2X1 NOR2X1_48 ( .A(_15_), .B(_372_), .Y(_373_) );
NAND2X1 NAND2X1_60 ( .A(dw04_cs), .B(_368_), .Y(_375_) );
AND2X2 AND2X2_11 ( .A(_368_), .B(dw0c_cs), .Y(_377_) );
NAND2X1 NAND2X1_61 ( .A(internal_counter_0_), .B(_377_), .Y(_378_) );
OAI21X1 OAI21X1_90 ( .A(_373__bF_buf2), .B(_378_), .C(_375_), .Y(_379_) );
AOI21X1 AOI21X1_25 ( .A(reg_08_data_0_), .B(_373__bF_buf2), .C(_379_), .Y(_380_) );
OAI21X1 OAI21X1_91 ( .A(reg_ito), .B(_375_), .C(_370_), .Y(_381_) );
OAI22X1 OAI22X1_15 ( .A(_364_), .B(_370_), .C(_381_), .D(_380_), .Y(_426__0_) );
INVX1 INVX1_50 ( .A(reg_run), .Y(_382_) );
NOR2X1 NOR2X1_49 ( .A(dw08_cs), .B(_98_), .Y(_383_) );
INVX1 INVX1_51 ( .A(_373__bF_buf2), .Y(_385_) );
OAI21X1 OAI21X1_92 ( .A(_100_), .B(_385_), .C(_375_), .Y(_386_) );
AOI21X1 AOI21X1_26 ( .A(_377_), .B(_383_), .C(_386_), .Y(_387_) );
OAI21X1 OAI21X1_93 ( .A(reg_cont), .B(_375_), .C(_370_), .Y(_388_) );
OAI22X1 OAI22X1_16 ( .A(_382_), .B(_370_), .C(_388_), .D(_387_), .Y(_426__1_) );
OAI21X1 OAI21X1_94 ( .A(dw04_cs), .B(dw00_cs), .C(_368_), .Y(_390_) );
INVX4 INVX4_6 ( .A(_390_), .Y(_391_) );
AND2X2 AND2X2_12 ( .A(_377_), .B(_15_), .Y(_392_) );
AOI22X1 AOI22X1_18 ( .A(reg_08_data_2_), .B(_373__bF_buf1), .C(internal_counter_2_), .D(_392_), .Y(_393_) );
NOR2X1 NOR2X1_50 ( .A(_391_), .B(_393_), .Y(_426__2_) );
AOI22X1 AOI22X1_19 ( .A(reg_08_data_3_), .B(_373__bF_buf0), .C(internal_counter_3_), .D(_392_), .Y(_394_) );
NOR2X1 NOR2X1_51 ( .A(_391_), .B(_394_), .Y(_426__3_) );
AOI22X1 AOI22X1_20 ( .A(reg_08_data_4_), .B(_373__bF_buf3), .C(internal_counter_4_), .D(_392_), .Y(_395_) );
NOR2X1 NOR2X1_52 ( .A(_391_), .B(_395_), .Y(_426__4_) );
AOI22X1 AOI22X1_21 ( .A(reg_08_data_5_), .B(_373__bF_buf1), .C(internal_counter_5_), .D(_392_), .Y(_396_) );
NOR2X1 NOR2X1_53 ( .A(_391_), .B(_396_), .Y(_426__5_) );
AOI22X1 AOI22X1_22 ( .A(reg_08_data_6_), .B(_373__bF_buf1), .C(internal_counter_6_), .D(_392_), .Y(_397_) );
NOR2X1 NOR2X1_54 ( .A(_391_), .B(_397_), .Y(_426__6_) );
AOI22X1 AOI22X1_23 ( .A(reg_08_data_7_), .B(_373__bF_buf1), .C(internal_counter_7_), .D(_392_), .Y(_398_) );
NOR2X1 NOR2X1_55 ( .A(_391_), .B(_398_), .Y(_426__7_) );
AOI22X1 AOI22X1_24 ( .A(reg_08_data_8_), .B(_373__bF_buf3), .C(internal_counter_8_), .D(_392_), .Y(_399_) );
NOR2X1 NOR2X1_56 ( .A(_391_), .B(_399_), .Y(_426__8_) );
AOI22X1 AOI22X1_25 ( .A(reg_08_data_9_), .B(_373__bF_buf3), .C(internal_counter_9_), .D(_392_), .Y(_400_) );
NOR2X1 NOR2X1_57 ( .A(_391_), .B(_400_), .Y(_426__9_) );
AOI22X1 AOI22X1_26 ( .A(reg_08_data_10_), .B(_373__bF_buf3), .C(internal_counter_10_), .D(_392_), .Y(_401_) );
NOR2X1 NOR2X1_58 ( .A(_391_), .B(_401_), .Y(_426__10_) );
AOI22X1 AOI22X1_27 ( .A(reg_08_data_11_), .B(_373__bF_buf3), .C(internal_counter_11_), .D(_392_), .Y(_402_) );
NOR2X1 NOR2X1_59 ( .A(_391_), .B(_402_), .Y(_426__11_) );
AOI22X1 AOI22X1_28 ( .A(reg_08_data_12_), .B(_373__bF_buf0), .C(internal_counter_12_), .D(_392_), .Y(_403_) );
NOR2X1 NOR2X1_60 ( .A(_391_), .B(_403_), .Y(_426__12_) );
AOI22X1 AOI22X1_29 ( .A(reg_08_data_13_), .B(_373__bF_buf0), .C(internal_counter_13_), .D(_392_), .Y(_404_) );
NOR2X1 NOR2X1_61 ( .A(_391_), .B(_404_), .Y(_426__13_) );
AOI22X1 AOI22X1_30 ( .A(reg_08_data_14_), .B(_373__bF_buf0), .C(internal_counter_14_), .D(_392_), .Y(_405_) );
NOR2X1 NOR2X1_62 ( .A(_391_), .B(_405_), .Y(_426__14_) );
AOI22X1 AOI22X1_31 ( .A(reg_08_data_15_), .B(_373__bF_buf2), .C(internal_counter_15_), .D(_392_), .Y(_406_) );
NOR2X1 NOR2X1_63 ( .A(_391_), .B(_406_), .Y(_426__15_) );
OAI21X1 OAI21X1_95 ( .A(_82_), .B(_51__bF_buf5), .C(_61_), .Y(_6__0_) );
OAI21X1 OAI21X1_96 ( .A(_100_), .B(_51__bF_buf3), .C(_96_), .Y(_6__1_) );
OAI21X1 OAI21X1_97 ( .A(_135_), .B(_51__bF_buf3), .C(_113_), .Y(_6__2_) );
OAI21X1 OAI21X1_98 ( .A(_136_), .B(_51__bF_buf5), .C(_132_), .Y(_6__3_) );
OAI21X1 OAI21X1_99 ( .A(_151_), .B(_51__bF_buf4), .C(_149_), .Y(_6__4_) );
INVX1 INVX1_52 ( .A(reg_08_data_5_), .Y(_407_) );
OAI21X1 OAI21X1_100 ( .A(_407_), .B(_51__bF_buf4), .C(_176_), .Y(_363_) );
OAI21X1 OAI21X1_101 ( .A(_193_), .B(_51__bF_buf4), .C(_189_), .Y(_365_) );
OAI21X1 OAI21X1_102 ( .A(_209_), .B(_51__bF_buf2), .C(_207_), .Y(_367_) );
OAI21X1 OAI21X1_103 ( .A(_225_), .B(_51__bF_buf2), .C(_224_), .Y(_369_) );
OAI21X1 OAI21X1_104 ( .A(_241_), .B(_51__bF_buf0), .C(_240_), .Y(_371_) );
OAI21X1 OAI21X1_105 ( .A(_262_), .B(_51__bF_buf0), .C(_260_), .Y(_6__10_) );
INVX1 INVX1_53 ( .A(reg_08_data_11_), .Y(_408_) );
OAI21X1 OAI21X1_106 ( .A(_408_), .B(_51__bF_buf2), .C(_288_), .Y(_374_) );
OAI21X1 OAI21X1_107 ( .A(_292_), .B(_51__bF_buf1), .C(_301_), .Y(_376_) );
NAND2X1 NAND2X1_62 ( .A(_325_), .B(_319_), .Y(_6__13_) );
OAI21X1 OAI21X1_108 ( .A(_74_), .B(_51__bF_buf1), .C(_330_), .Y(_6__14_) );
OAI21X1 OAI21X1_109 ( .A(_75_), .B(_51__bF_buf1), .C(_354_), .Y(_6__15_) );
INVX1 INVX1_54 ( .A(dw04_cs), .Y(_409_) );
NOR2X1 NOR2X1_64 ( .A(_16_), .B(_409_), .Y(_410_) );
INVX2 INVX2_12 ( .A(_410_), .Y(_411_) );
OAI21X1 OAI21X1_110 ( .A(latch_s_data_3_), .B(_411_), .C(reg_stop), .Y(_412_) );
NOR2X1 NOR2X1_65 ( .A(latch_s_data_2_), .B(_411_), .Y(_413_) );
OAI21X1 OAI21X1_111 ( .A(reg_stop), .B(latch_s_data_3_), .C(_413_), .Y(_414_) );
NAND2X1 NAND2X1_63 ( .A(_412_), .B(_414_), .Y(_384_) );
OAI21X1 OAI21X1_112 ( .A(status_2_), .B(status_1_bF_buf0), .C(_40_), .Y(_415_) );
OAI21X1 OAI21X1_113 ( .A(reg_stop), .B(_12_), .C(_415_), .Y(_7_) );
INVX1 INVX1_55 ( .A(latch_s_data_0_), .Y(_416_) );
OAI21X1 OAI21X1_114 ( .A(_16_), .B(_409_), .C(reg_ito), .Y(_417_) );
OAI21X1 OAI21X1_115 ( .A(_416_), .B(_411_), .C(_417_), .Y(_5__0_) );
NAND2X1 NAND2X1_64 ( .A(latch_s_data_1_), .B(_410_), .Y(_418_) );
OAI21X1 OAI21X1_116 ( .A(_47_), .B(_410_), .C(_418_), .Y(_389_) );
NAND3X1 NAND3X1_39 ( .A(reg_run), .B(reg_ito), .C(_41_), .Y(_419_) );
NOR2X1 NOR2X1_66 ( .A(latch_s_data_0_), .B(_16_), .Y(_420_) );
AOI22X1 AOI22X1_32 ( .A(dw00_cs), .B(_420_), .C(_364_), .D(_419_), .Y(_9_) );
INVX1 INVX1_56 ( .A(s_ack_dly), .Y(_421_) );
NOR2X1 NOR2X1_67 ( .A(s_ack_2dly), .B(_421_), .Y(_425_) );
NAND2X1 NAND2X1_65 ( .A(latch_s_data_2_), .B(_382_), .Y(_422_) );
NOR2X1 NOR2X1_68 ( .A(_422_), .B(_411_), .Y(_8_) );
INVX8 INVX8_1 ( .A(RST_I), .Y(_429_) );
BUFX2 BUFX2_8 ( .A(_undef), .Y(RSTREQ_O) );
BUFX2 BUFX2_9 ( .A(_425_), .Y(S_ACK_O) );
BUFX2 BUFX2_10 ( .A(_426__0_), .Y(S_DAT_O[0]) );
BUFX2 BUFX2_11 ( .A(_426__1_), .Y(S_DAT_O[1]) );
BUFX2 BUFX2_12 ( .A(_426__2_), .Y(S_DAT_O[2]) );
BUFX2 BUFX2_13 ( .A(_426__3_), .Y(S_DAT_O[3]) );
BUFX2 BUFX2_14 ( .A(_426__4_), .Y(S_DAT_O[4]) );
BUFX2 BUFX2_15 ( .A(_426__5_), .Y(S_DAT_O[5]) );
BUFX2 BUFX2_16 ( .A(_426__6_), .Y(S_DAT_O[6]) );
BUFX2 BUFX2_17 ( .A(_426__7_), .Y(S_DAT_O[7]) );
BUFX2 BUFX2_18 ( .A(_426__8_), .Y(S_DAT_O[8]) );
BUFX2 BUFX2_19 ( .A(_426__9_), .Y(S_DAT_O[9]) );
BUFX2 BUFX2_20 ( .A(_426__10_), .Y(S_DAT_O[10]) );
BUFX2 BUFX2_21 ( .A(_426__11_), .Y(S_DAT_O[11]) );
BUFX2 BUFX2_22 ( .A(_426__12_), .Y(S_DAT_O[12]) );
BUFX2 BUFX2_23 ( .A(_426__13_), .Y(S_DAT_O[13]) );
BUFX2 BUFX2_24 ( .A(_426__14_), .Y(S_DAT_O[14]) );
BUFX2 BUFX2_25 ( .A(_426__15_), .Y(S_DAT_O[15]) );
BUFX2 BUFX2_26 ( .A(gnd), .Y(S_DAT_O[16]) );
BUFX2 BUFX2_27 ( .A(gnd), .Y(S_DAT_O[17]) );
BUFX2 BUFX2_28 ( .A(gnd), .Y(S_DAT_O[18]) );
BUFX2 BUFX2_29 ( .A(gnd), .Y(S_DAT_O[19]) );
BUFX2 BUFX2_30 ( .A(gnd), .Y(S_DAT_O[20]) );
BUFX2 BUFX2_31 ( .A(gnd), .Y(S_DAT_O[21]) );
BUFX2 BUFX2_32 ( .A(gnd), .Y(S_DAT_O[22]) );
BUFX2 BUFX2_33 ( .A(gnd), .Y(S_DAT_O[23]) );
BUFX2 BUFX2_34 ( .A(gnd), .Y(S_DAT_O[24]) );
BUFX2 BUFX2_35 ( .A(gnd), .Y(S_DAT_O[25]) );
BUFX2 BUFX2_36 ( .A(gnd), .Y(S_DAT_O[26]) );
BUFX2 BUFX2_37 ( .A(gnd), .Y(S_DAT_O[27]) );
BUFX2 BUFX2_38 ( .A(gnd), .Y(S_DAT_O[28]) );
BUFX2 BUFX2_39 ( .A(gnd), .Y(S_DAT_O[29]) );
BUFX2 BUFX2_40 ( .A(gnd), .Y(S_DAT_O[30]) );
BUFX2 BUFX2_41 ( .A(gnd), .Y(S_DAT_O[31]) );
BUFX2 BUFX2_42 ( .A(gnd), .Y(S_ERR_O) );
BUFX2 BUFX2_43 ( .A(_427_), .Y(S_INT_O) );
BUFX2 BUFX2_44 ( .A(gnd), .Y(S_RTY_O) );
BUFX2 BUFX2_45 ( .A(_428_), .Y(TOPULSE_O) );
DFFSR DFFSR_1 ( .CLK(CLK_I_bF_buf4), .D(_424__0_), .Q(status_0_), .R(vdd), .S(_429__bF_buf5) );
DFFSR DFFSR_2 ( .CLK(CLK_I_bF_buf4), .D(_424__1_), .Q(status_1_), .R(_429__bF_buf7), .S(vdd) );
DFFSR DFFSR_3 ( .CLK(CLK_I_bF_buf0), .D(_424__2_), .Q(status_2_), .R(_429__bF_buf0), .S(vdd) );
DFFSR DFFSR_4 ( .CLK(CLK_I_bF_buf6), .D(_423_), .Q(_428_), .R(_429__bF_buf6), .S(vdd) );
DFFSR DFFSR_5 ( .CLK(CLK_I_bF_buf6), .D(_6__0_), .Q(reg_08_data_0_), .R(_429__bF_buf0), .S(vdd) );
DFFSR DFFSR_6 ( .CLK(CLK_I_bF_buf7), .D(_6__1_), .Q(reg_08_data_1_), .R(_429__bF_buf4), .S(vdd) );
DFFSR DFFSR_7 ( .CLK(CLK_I_bF_buf7), .D(_6__2_), .Q(reg_08_data_2_), .R(vdd), .S(_429__bF_buf2) );
DFFSR DFFSR_8 ( .CLK(CLK_I_bF_buf0), .D(_6__3_), .Q(reg_08_data_3_), .R(_429__bF_buf5), .S(vdd) );
DFFSR DFFSR_9 ( .CLK(CLK_I_bF_buf4), .D(_6__4_), .Q(reg_08_data_4_), .R(vdd), .S(_429__bF_buf7) );
DFFSR DFFSR_10 ( .CLK(CLK_I_bF_buf4), .D(_363_), .Q(reg_08_data_5_), .R(_429__bF_buf7), .S(vdd) );
DFFSR DFFSR_11 ( .CLK(CLK_I_bF_buf1), .D(_365_), .Q(reg_08_data_6_), .R(_429__bF_buf3), .S(vdd) );
DFFSR DFFSR_12 ( .CLK(CLK_I_bF_buf1), .D(_367_), .Q(reg_08_data_7_), .R(_429__bF_buf3), .S(vdd) );
DFFSR DFFSR_13 ( .CLK(CLK_I_bF_buf2), .D(_369_), .Q(reg_08_data_8_), .R(_429__bF_buf7), .S(vdd) );
DFFSR DFFSR_14 ( .CLK(CLK_I_bF_buf5), .D(_371_), .Q(reg_08_data_9_), .R(_429__bF_buf1), .S(vdd) );
DFFSR DFFSR_15 ( .CLK(CLK_I_bF_buf2), .D(_6__10_), .Q(reg_08_data_10_), .R(_429__bF_buf1), .S(vdd) );
DFFSR DFFSR_16 ( .CLK(CLK_I_bF_buf1), .D(_374_), .Q(reg_08_data_11_), .R(_429__bF_buf3), .S(vdd) );
DFFSR DFFSR_17 ( .CLK(CLK_I_bF_buf5), .D(_376_), .Q(reg_08_data_12_), .R(_429__bF_buf5), .S(vdd) );
DFFSR DFFSR_18 ( .CLK(CLK_I_bF_buf5), .D(_6__13_), .Q(reg_08_data_13_), .R(_429__bF_buf5), .S(vdd) );
DFFSR DFFSR_19 ( .CLK(CLK_I_bF_buf0), .D(_6__14_), .Q(reg_08_data_14_), .R(_429__bF_buf0), .S(vdd) );
DFFSR DFFSR_20 ( .CLK(CLK_I_bF_buf0), .D(_6__15_), .Q(reg_08_data_15_), .R(_429__bF_buf5), .S(vdd) );
DFFSR DFFSR_21 ( .CLK(CLK_I_bF_buf6), .D(_384_), .Q(reg_stop), .R(_429__bF_buf6), .S(vdd) );
DFFSR DFFSR_22 ( .CLK(CLK_I_bF_buf0), .D(_7_), .Q(reg_run), .R(_429__bF_buf0), .S(vdd) );
DFFSR DFFSR_23 ( .CLK(CLK_I_bF_buf3), .D(_14_), .Q(internal_counter_0_), .R(_429__bF_buf4), .S(vdd) );
DFFSR DFFSR_24 ( .CLK(CLK_I_bF_buf7), .D(_31_), .Q(internal_counter_1_), .R(_429__bF_buf2), .S(vdd) );
DFFSR DFFSR_25 ( .CLK(CLK_I_bF_buf7), .D(_48_), .Q(internal_counter_2_), .R(_429__bF_buf2), .S(vdd) );
DFFSR DFFSR_26 ( .CLK(CLK_I_bF_buf3), .D(_60_), .Q(internal_counter_3_), .R(_429__bF_buf6), .S(vdd) );
DFFSR DFFSR_27 ( .CLK(CLK_I_bF_buf4), .D(_81_), .Q(internal_counter_4_), .R(_429__bF_buf7), .S(vdd) );
DFFSR DFFSR_28 ( .CLK(CLK_I_bF_buf2), .D(_99_), .Q(internal_counter_5_), .R(_429__bF_buf7), .S(vdd) );
DFFSR DFFSR_29 ( .CLK(CLK_I_bF_buf4), .D(_120_), .Q(internal_counter_6_), .R(_429__bF_buf7), .S(vdd) );
DFFSR DFFSR_30 ( .CLK(CLK_I_bF_buf1), .D(_138_), .Q(internal_counter_7_), .R(_429__bF_buf3), .S(vdd) );
DFFSR DFFSR_31 ( .CLK(CLK_I_bF_buf2), .D(_161_), .Q(internal_counter_8_), .R(_429__bF_buf1), .S(vdd) );
DFFSR DFFSR_32 ( .CLK(CLK_I_bF_buf2), .D(_179_), .Q(internal_counter_9_), .R(_429__bF_buf7), .S(vdd) );
DFFSR DFFSR_33 ( .CLK(CLK_I_bF_buf2), .D(_204_), .Q(internal_counter_10_), .R(_429__bF_buf1), .S(vdd) );
DFFSR DFFSR_34 ( .CLK(CLK_I_bF_buf2), .D(_222_), .Q(internal_counter_11_), .R(_429__bF_buf7), .S(vdd) );
DFFSR DFFSR_35 ( .CLK(CLK_I_bF_buf5), .D(_243_), .Q(internal_counter_12_), .R(_429__bF_buf5), .S(vdd) );
DFFSR DFFSR_36 ( .CLK(CLK_I_bF_buf5), .D(_261_), .Q(internal_counter_13_), .R(_429__bF_buf1), .S(vdd) );
DFFSR DFFSR_37 ( .CLK(CLK_I_bF_buf0), .D(_4__14_), .Q(internal_counter_14_), .R(_429__bF_buf0), .S(vdd) );
DFFSR DFFSR_38 ( .CLK(CLK_I_bF_buf4), .D(_4__15_), .Q(internal_counter_15_), .R(_429__bF_buf2), .S(vdd) );
DFFSR DFFSR_39 ( .CLK(CLK_I_bF_buf7), .D(s_ack_pre), .Q(s_ack_dly), .R(_429__bF_buf2), .S(vdd) );
DFFSR DFFSR_40 ( .CLK(CLK_I_bF_buf7), .D(s_ack_dly), .Q(s_ack_2dly), .R(_429__bF_buf2), .S(vdd) );
DFFSR DFFSR_41 ( .CLK(CLK_I_bF_buf7), .D(_11_), .Q(s_ack_pre), .R(_429__bF_buf4), .S(vdd) );
DFFSR DFFSR_42 ( .CLK(CLK_I_bF_buf6), .D(_5__0_), .Q(reg_ito), .R(_429__bF_buf6), .S(vdd) );
DFFSR DFFSR_43 ( .CLK(CLK_I_bF_buf3), .D(_389_), .Q(reg_cont), .R(_429__bF_buf6), .S(vdd) );
DFFSR DFFSR_44 ( .CLK(CLK_I_bF_buf6), .D(_8_), .Q(reg_start), .R(_429__bF_buf0), .S(vdd) );
DFFSR DFFSR_45 ( .CLK(CLK_I_bF_buf3), .D(_9_), .Q(_427_), .R(_429__bF_buf6), .S(vdd) );
DFFSR DFFSR_46 ( .CLK(CLK_I_bF_buf6), .D(_10_), .Q(reg_wr), .R(_429__bF_buf6), .S(vdd) );
DFFSR DFFSR_47 ( .CLK(CLK_I_bF_buf3), .D(_0_), .Q(dw00_cs), .R(_429__bF_buf4), .S(vdd) );
DFFSR DFFSR_48 ( .CLK(CLK_I_bF_buf3), .D(_1_), .Q(dw04_cs), .R(_429__bF_buf4), .S(vdd) );
DFFSR DFFSR_49 ( .CLK(CLK_I_bF_buf3), .D(_2_), .Q(dw08_cs), .R(_429__bF_buf4), .S(vdd) );
DFFSR DFFSR_50 ( .CLK(CLK_I_bF_buf3), .D(_3_), .Q(dw0c_cs), .R(_429__bF_buf4), .S(vdd) );
DFFSR DFFSR_51 ( .CLK(CLK_I_bF_buf7), .D(S_DAT_I[0]), .Q(latch_s_data_0_), .R(_429__bF_buf4), .S(vdd) );
DFFSR DFFSR_52 ( .CLK(CLK_I_bF_buf6), .D(S_DAT_I[1]), .Q(latch_s_data_1_), .R(_429__bF_buf0), .S(vdd) );
DFFSR DFFSR_53 ( .CLK(CLK_I_bF_buf6), .D(S_DAT_I[2]), .Q(latch_s_data_2_), .R(_429__bF_buf6), .S(vdd) );
DFFSR DFFSR_54 ( .CLK(CLK_I_bF_buf6), .D(S_DAT_I[3]), .Q(latch_s_data_3_), .R(_429__bF_buf6), .S(vdd) );
DFFSR DFFSR_55 ( .CLK(CLK_I_bF_buf1), .D(S_DAT_I[4]), .Q(latch_s_data_4_), .R(_429__bF_buf3), .S(vdd) );
DFFSR DFFSR_56 ( .CLK(CLK_I_bF_buf0), .D(S_DAT_I[5]), .Q(latch_s_data_5_), .R(_429__bF_buf0), .S(vdd) );
DFFSR DFFSR_57 ( .CLK(CLK_I_bF_buf1), .D(S_DAT_I[6]), .Q(latch_s_data_6_), .R(_429__bF_buf3), .S(vdd) );
DFFSR DFFSR_58 ( .CLK(CLK_I_bF_buf1), .D(S_DAT_I[7]), .Q(latch_s_data_7_), .R(_429__bF_buf3), .S(vdd) );
DFFSR DFFSR_59 ( .CLK(CLK_I_bF_buf1), .D(S_DAT_I[8]), .Q(latch_s_data_8_), .R(_429__bF_buf3), .S(vdd) );
DFFSR DFFSR_60 ( .CLK(CLK_I_bF_buf5), .D(S_DAT_I[9]), .Q(latch_s_data_9_), .R(_429__bF_buf5), .S(vdd) );
DFFSR DFFSR_61 ( .CLK(CLK_I_bF_buf2), .D(S_DAT_I[10]), .Q(latch_s_data_10_), .R(_429__bF_buf1), .S(vdd) );
DFFSR DFFSR_62 ( .CLK(CLK_I_bF_buf4), .D(S_DAT_I[11]), .Q(latch_s_data_11_), .R(_429__bF_buf2), .S(vdd) );
DFFSR DFFSR_63 ( .CLK(CLK_I_bF_buf5), .D(S_DAT_I[12]), .Q(latch_s_data_12_), .R(_429__bF_buf1), .S(vdd) );
DFFSR DFFSR_64 ( .CLK(CLK_I_bF_buf5), .D(S_DAT_I[13]), .Q(latch_s_data_13_), .R(_429__bF_buf1), .S(vdd) );
DFFSR DFFSR_65 ( .CLK(CLK_I_bF_buf0), .D(S_DAT_I[14]), .Q(latch_s_data_14_), .R(_429__bF_buf5), .S(vdd) );
DFFSR DFFSR_66 ( .CLK(CLK_I_bF_buf7), .D(S_DAT_I[15]), .Q(latch_s_data_15_), .R(_429__bF_buf2), .S(vdd) );
endmodule
